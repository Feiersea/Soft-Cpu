module Register (
    input wire enable;
    input wire clk;
    input wire reg_in1;
    output reg reg_out1;

);